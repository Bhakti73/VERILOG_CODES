timescale 1ns / 1ps

module gates(
input a,
output y
    );
    
    assign y = ~a;
    
endmodule